//Test Bench:
// THIS IS A TEST BENCH FOR SIMPLE UN PIPELINED FLOATING POINT ADDER
/*
SET of INPUTS and expected outputs:
1.
    100=01000010110010000000000000000000
    200=01000011010010000000000000000000
    300=01000011100101100000000000000000

2.
    100=01000010110010000000000000000000
   -50= 11000010010010000000000000000000
    50= 01000010010010000000000000000000
3. 
    -53= 11000010010101000000000000000000
    -35=11000010000011000000000000000000
    -88=11000010101100000000000000000000
4.
    -300=11000011100101100000000000000000
    -99=11000010110001100000000000000000
    -399=11000011110001111000000000000000
5.
    0=00000000000000000000000000000000
    
6. 
    0-171= 
    -171=11000011001010110000000000000000
*/

module tb_unfp_40 ();
reg  [31:0]  a,b;
wire [31:0] r;
reg clk, rst;
unfp_40 t(a,b,r,rst,clk);
initial begin
clk = 0;
rst = 0;
#2;
rst = 1;
#2;
rst = 0;
end
initial forever #5 clk = ~clk;
initial begin
// 1st input:
#10
a= 32'b01000010110010000000000000000000;
b= 32'b01000011010010000000000000000000; 
// 2nd input:
#10
$display("result is : %b",  r);
a= 32'b01000010110010000000000000000000;
b= 32'b11000010010010000000000000000000; 
// 3rd input:
#10
$display("result is : %b",  r);
a= 32'b11000010010101000000000000000000;
b= 32'b11000010000011000000000000000000; 
//4 input
#10
$display("result is : %b",  r);
a= 32'b11000011100101100000000000000000;
b= 32'b11000010110001100000000000000000; 
//5 input
#10
$display("result is : %b",  r);
a= 32'b00000000000000000000000000000000;
b= 32'b00000000000000000000000000000000; 
//6 input
#10
$display("result is : %b",  r);
a= 32'b00000000000000000000000000000000;
b= 32'b11000011001010110000000000000000; 
#10
$display("result is : %b",  r);
$finish;
end
initial begin 
$dumpfile ("1a.vcd");
$dumpvars (0,tb_unfp_40);
end
endmodule
